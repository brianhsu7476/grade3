module Add(a, b, c);
input signed[31:0]a, b;
output signed[31:0]c;
assign c=a+b;
endmodule
